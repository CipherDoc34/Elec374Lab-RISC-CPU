library verilog;
use verilog.vl_types.all;
entity datapath_tb is
    generic(
        Default         : integer := 0;
        Reg_load1a      : integer := 1;
        Reg_load1b      : integer := 2;
        Reg_load2a      : integer := 3;
        Reg_load2b      : integer := 4;
        Reg_load3a      : integer := 5;
        Reg_load3b      : integer := 6;
        Reg_load4a      : integer := 7;
        Reg_load4b      : integer := 8;
        Reg_load5a      : integer := 9;
        Reg_load5b      : integer := 10;
        Reg_load6a      : integer := 11;
        Reg_load6b      : integer := 12;
        Reg_load7a      : integer := 13;
        Reg_load7b      : integer := 14;
        ANDT0           : integer := 15;
        ANDT1           : integer := 16;
        ANDT2           : integer := 17;
        ANDT3           : integer := 18;
        ANDT4           : integer := 19;
        ANDT5           : integer := 20;
        ADDT0           : integer := 21;
        ADDT1           : integer := 22;
        ADDT2           : integer := 23;
        ADDT3           : integer := 24;
        ADDT4           : integer := 25;
        ADDT5           : integer := 26;
        SUBT0           : integer := 27;
        SUBT1           : integer := 28;
        SUBT2           : integer := 29;
        SUBT3           : integer := 30;
        SUBT4           : integer := 31;
        SUBT5           : integer := 32;
        MULT0           : integer := 33;
        MULT1           : integer := 34;
        MULT2           : integer := 35;
        MULT3           : integer := 36;
        MULT4           : integer := 37;
        MULT5           : integer := 38;
        MULT6           : integer := 39;
        DIVT0           : integer := 40;
        DIVT1           : integer := 41;
        DIVT2           : integer := 42;
        DIVT3           : integer := 43;
        DIVT4           : integer := 44;
        DIVT5           : integer := 45;
        DIVT6           : integer := 46;
        SHRT0           : integer := 47;
        SHRT1           : integer := 48;
        SHRT2           : integer := 49;
        SHRT3           : integer := 50;
        SHRT4           : integer := 51;
        SHRT5           : integer := 52;
        SHRAT0          : integer := 53;
        SHRAT1          : integer := 54;
        SHRAT2          : integer := 55;
        SHRAT3          : integer := 56;
        SHRAT4          : integer := 57;
        SHRAT5          : integer := 58;
        SHLT0           : integer := 59;
        SHLT1           : integer := 60;
        SHLT2           : integer := 61;
        SHLT3           : integer := 62;
        SHLT4           : integer := 63;
        SHLT5           : integer := 64;
        RORT0           : integer := 65;
        RORT1           : integer := 66;
        RORT2           : integer := 67;
        RORT3           : integer := 68;
        RORT4           : integer := 69;
        RORT5           : integer := 70;
        ROLT0           : integer := 71;
        ROLT1           : integer := 72;
        ROLT2           : integer := 73;
        ROLT3           : integer := 74;
        ROLT4           : integer := 75;
        ROLT5           : integer := 76;
        NEGT0           : integer := 77;
        NEGT1           : integer := 78;
        NEGT2           : integer := 79;
        NEGT3           : integer := 80;
        NEGT4           : integer := 81;
        NEGT5           : integer := 82;
        NOTT0           : integer := 83;
        NOTT1           : integer := 84;
        NOTT2           : integer := 85;
        NOTT3           : integer := 86;
        NOTT4           : integer := 87;
        NOTT5           : integer := 88
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of Default : constant is 1;
    attribute mti_svvh_generic_type of Reg_load1a : constant is 1;
    attribute mti_svvh_generic_type of Reg_load1b : constant is 1;
    attribute mti_svvh_generic_type of Reg_load2a : constant is 1;
    attribute mti_svvh_generic_type of Reg_load2b : constant is 1;
    attribute mti_svvh_generic_type of Reg_load3a : constant is 1;
    attribute mti_svvh_generic_type of Reg_load3b : constant is 1;
    attribute mti_svvh_generic_type of Reg_load4a : constant is 1;
    attribute mti_svvh_generic_type of Reg_load4b : constant is 1;
    attribute mti_svvh_generic_type of Reg_load5a : constant is 1;
    attribute mti_svvh_generic_type of Reg_load5b : constant is 1;
    attribute mti_svvh_generic_type of Reg_load6a : constant is 1;
    attribute mti_svvh_generic_type of Reg_load6b : constant is 1;
    attribute mti_svvh_generic_type of Reg_load7a : constant is 1;
    attribute mti_svvh_generic_type of Reg_load7b : constant is 1;
    attribute mti_svvh_generic_type of ANDT0 : constant is 1;
    attribute mti_svvh_generic_type of ANDT1 : constant is 1;
    attribute mti_svvh_generic_type of ANDT2 : constant is 1;
    attribute mti_svvh_generic_type of ANDT3 : constant is 1;
    attribute mti_svvh_generic_type of ANDT4 : constant is 1;
    attribute mti_svvh_generic_type of ANDT5 : constant is 1;
    attribute mti_svvh_generic_type of ADDT0 : constant is 1;
    attribute mti_svvh_generic_type of ADDT1 : constant is 1;
    attribute mti_svvh_generic_type of ADDT2 : constant is 1;
    attribute mti_svvh_generic_type of ADDT3 : constant is 1;
    attribute mti_svvh_generic_type of ADDT4 : constant is 1;
    attribute mti_svvh_generic_type of ADDT5 : constant is 1;
    attribute mti_svvh_generic_type of SUBT0 : constant is 1;
    attribute mti_svvh_generic_type of SUBT1 : constant is 1;
    attribute mti_svvh_generic_type of SUBT2 : constant is 1;
    attribute mti_svvh_generic_type of SUBT3 : constant is 1;
    attribute mti_svvh_generic_type of SUBT4 : constant is 1;
    attribute mti_svvh_generic_type of SUBT5 : constant is 1;
    attribute mti_svvh_generic_type of MULT0 : constant is 1;
    attribute mti_svvh_generic_type of MULT1 : constant is 1;
    attribute mti_svvh_generic_type of MULT2 : constant is 1;
    attribute mti_svvh_generic_type of MULT3 : constant is 1;
    attribute mti_svvh_generic_type of MULT4 : constant is 1;
    attribute mti_svvh_generic_type of MULT5 : constant is 1;
    attribute mti_svvh_generic_type of MULT6 : constant is 1;
    attribute mti_svvh_generic_type of DIVT0 : constant is 1;
    attribute mti_svvh_generic_type of DIVT1 : constant is 1;
    attribute mti_svvh_generic_type of DIVT2 : constant is 1;
    attribute mti_svvh_generic_type of DIVT3 : constant is 1;
    attribute mti_svvh_generic_type of DIVT4 : constant is 1;
    attribute mti_svvh_generic_type of DIVT5 : constant is 1;
    attribute mti_svvh_generic_type of DIVT6 : constant is 1;
    attribute mti_svvh_generic_type of SHRT0 : constant is 1;
    attribute mti_svvh_generic_type of SHRT1 : constant is 1;
    attribute mti_svvh_generic_type of SHRT2 : constant is 1;
    attribute mti_svvh_generic_type of SHRT3 : constant is 1;
    attribute mti_svvh_generic_type of SHRT4 : constant is 1;
    attribute mti_svvh_generic_type of SHRT5 : constant is 1;
    attribute mti_svvh_generic_type of SHRAT0 : constant is 1;
    attribute mti_svvh_generic_type of SHRAT1 : constant is 1;
    attribute mti_svvh_generic_type of SHRAT2 : constant is 1;
    attribute mti_svvh_generic_type of SHRAT3 : constant is 1;
    attribute mti_svvh_generic_type of SHRAT4 : constant is 1;
    attribute mti_svvh_generic_type of SHRAT5 : constant is 1;
    attribute mti_svvh_generic_type of SHLT0 : constant is 1;
    attribute mti_svvh_generic_type of SHLT1 : constant is 1;
    attribute mti_svvh_generic_type of SHLT2 : constant is 1;
    attribute mti_svvh_generic_type of SHLT3 : constant is 1;
    attribute mti_svvh_generic_type of SHLT4 : constant is 1;
    attribute mti_svvh_generic_type of SHLT5 : constant is 1;
    attribute mti_svvh_generic_type of RORT0 : constant is 1;
    attribute mti_svvh_generic_type of RORT1 : constant is 1;
    attribute mti_svvh_generic_type of RORT2 : constant is 1;
    attribute mti_svvh_generic_type of RORT3 : constant is 1;
    attribute mti_svvh_generic_type of RORT4 : constant is 1;
    attribute mti_svvh_generic_type of RORT5 : constant is 1;
    attribute mti_svvh_generic_type of ROLT0 : constant is 1;
    attribute mti_svvh_generic_type of ROLT1 : constant is 1;
    attribute mti_svvh_generic_type of ROLT2 : constant is 1;
    attribute mti_svvh_generic_type of ROLT3 : constant is 1;
    attribute mti_svvh_generic_type of ROLT4 : constant is 1;
    attribute mti_svvh_generic_type of ROLT5 : constant is 1;
    attribute mti_svvh_generic_type of NEGT0 : constant is 1;
    attribute mti_svvh_generic_type of NEGT1 : constant is 1;
    attribute mti_svvh_generic_type of NEGT2 : constant is 1;
    attribute mti_svvh_generic_type of NEGT3 : constant is 1;
    attribute mti_svvh_generic_type of NEGT4 : constant is 1;
    attribute mti_svvh_generic_type of NEGT5 : constant is 1;
    attribute mti_svvh_generic_type of NOTT0 : constant is 1;
    attribute mti_svvh_generic_type of NOTT1 : constant is 1;
    attribute mti_svvh_generic_type of NOTT2 : constant is 1;
    attribute mti_svvh_generic_type of NOTT3 : constant is 1;
    attribute mti_svvh_generic_type of NOTT4 : constant is 1;
    attribute mti_svvh_generic_type of NOTT5 : constant is 1;
end datapath_tb;
