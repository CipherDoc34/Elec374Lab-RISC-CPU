library verilog;
use verilog.vl_types.all;
entity \Bus\ is
    port(
        BusMuxInR0      : in     vl_logic_vector(31 downto 0);
        BusMuxInR1      : in     vl_logic_vector(31 downto 0);
        BusMuxInR2      : in     vl_logic_vector(31 downto 0);
        BusMuxInR3      : in     vl_logic_vector(31 downto 0);
        BusMuxInR4      : in     vl_logic_vector(31 downto 0);
        BusMuxInR5      : in     vl_logic_vector(31 downto 0);
        BusMuxInR6      : in     vl_logic_vector(31 downto 0);
        BusMuxInR7      : in     vl_logic_vector(31 downto 0);
        BusMuxInR8      : in     vl_logic_vector(31 downto 0);
        BusMuxInR9      : in     vl_logic_vector(31 downto 0);
        BusMuxInR10     : in     vl_logic_vector(31 downto 0);
        BusMuxInR11     : in     vl_logic_vector(31 downto 0);
        BusMuxInR12     : in     vl_logic_vector(31 downto 0);
        BusMuxInR13     : in     vl_logic_vector(31 downto 0);
        BusMuxInR14     : in     vl_logic_vector(31 downto 0);
        BusMuxInR15     : in     vl_logic_vector(31 downto 0);
        BusMuxInHI      : in     vl_logic_vector(31 downto 0);
        BusMuxInLO      : in     vl_logic_vector(31 downto 0);
        BusMuxInZHI     : in     vl_logic_vector(31 downto 0);
        BusMuxInZLO     : in     vl_logic_vector(31 downto 0);
        BusMuxInZMux    : in     vl_logic_vector(31 downto 0);
        BusMuxInPC      : in     vl_logic_vector(31 downto 0);
        BusMuxInMDR     : in     vl_logic_vector(31 downto 0);
        BusMuxInPortIn  : in     vl_logic_vector(31 downto 0);
        BusMuxInCSign   : in     vl_logic_vector(31 downto 0);
        R0out           : in     vl_logic;
        R1out           : in     vl_logic;
        R2out           : in     vl_logic;
        R3out           : in     vl_logic;
        R4out           : in     vl_logic;
        R5out           : in     vl_logic;
        R6out           : in     vl_logic;
        R7out           : in     vl_logic;
        R8out           : in     vl_logic;
        R9out           : in     vl_logic;
        R10out          : in     vl_logic;
        R11out          : in     vl_logic;
        R12out          : in     vl_logic;
        R13out          : in     vl_logic;
        R14out          : in     vl_logic;
        R15out          : in     vl_logic;
        HIout           : in     vl_logic;
        LOout           : in     vl_logic;
        ZHIout          : in     vl_logic;
        ZLOout          : in     vl_logic;
        ZMuxOut         : in     vl_logic;
        PCout           : in     vl_logic;
        MDRout          : in     vl_logic;
        PortInout       : in     vl_logic;
        CSignout        : in     vl_logic;
        S0              : out    vl_logic;
        S1              : out    vl_logic;
        S2              : out    vl_logic;
        S3              : out    vl_logic;
        S4              : out    vl_logic;
        BusMuxOut       : out    vl_logic_vector(31 downto 0)
    );
end \Bus\;
